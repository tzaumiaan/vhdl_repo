library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
library std;
use std.textio.all;

entity tb is
end entity tb;

architecture rtl of tb is
begin
end architecture rtl;
